`timescale 1ns / 1ps
`include "CPU_Param.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:00:54 11/22/2020 
// Design Name: 
// Module Name:    ID 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ID(
    input wire [31:0] Instr,
    input wire [31:0] PC,
    input wire [31:0] PC_4,
    input wire clk,
    input wire reset,
	input wire RegWrite,
	input wire [31:0] WData,
	input wire [31:0] WritePC,
	input wire [4:0] RegWriteAddr_Mem_to_WB,
    output reg [4:0] Rs_ID_to_EX,
    output reg [4:0] Rt_ID_to_EX,
    output reg [4:0] RegWriteAddr_ID_to_EX, //��ָ����Rd�����ǵ�ǰָ����ʵ����д���GPR��ַ
    output reg [4:0] Shamt_ID_to_EX,
    output reg [31:0] imm32_ID_to_EX,
	output reg [59:0] InstrType_ID_to_EX,
	output reg [31:0] RsData_ID_to_EX,
	output reg [31:0] RtData_ID_to_EX,
    output reg [31:0] luiRes_ID_to_EX,
	output reg [31:0] PC_ID_to_EX,
	output wire branch,
    output wire jump,
    output wire [31:0] branch_addr32,
    output wire [31:0] jump_addr32
    );
	wire [31:0] RsData_wire, RtData_wire, imm32_wire;
	wire [25:0] imm26_wire;
	wire [15:0] imm16_wire;
	wire [4:0] Rs_wire, Rt_wire, Rd_wire, Shamt_wire;
	wire sign;
	wire [59:0] InstrType;
	
	//ת����ûд����ת��������д�ú����RsData_wire��RtData_wire��MUX
	//�Լ�T_use��T_new
	
	assign sign = (`ori || `sll) ? 0 : 1 ; //�������Ӧ��0��չ��ָ�����
	assign {Rs_wire, Rt_wire, Rd_wire, Shamt_wire} = Instr[25:6];
	assign imm26_wire = Instr[25:0];
	assign imm16_wire = `sll ? {11'd0, Shamt_wire} : Instr[15:0];
	
	
	InstrDecoder InstrDecoder(
	.Instr(Instr),
	.InstrType(InstrType));
	
	Extender Extender(
	.imm16(imm16_wire),
	.sign(sign),
	.imm32(imm32_wire));
	
	wire [4:0] WAddr_wire;
	wire [31:0] RData0_wire, RData1_wire, RData0_read;
	assign WAddr_wire = (`jal) ? 5'd31 :
	               (`ori || `lw || `lui) ? Rt_wire : Rd_wire;
	// Instructions write to GPR No.31 or Rt
	GRF GRF(
	.RAddr0(Rs_wire),
	.RAddr1(Rt_wire),
	.WAddr(RegWriteAddr_Mem_to_WB),
	.WriteData(WData),
	.WritePC(WritePC), //дָ���PC���ǵ�ǰPC
	.RegWrite(RegWrite),
	.clk(clk),
	.reset(reset),
	.RData0(RData0_read), //ԭʼ��������
	.RData1(RData1_wire));
	assign RData0_wire = (`sll) ? {27'd0, Shamt_wire} : RData0_read;
	//����sll����Rs����Shamt��Ϊsllv��ʣ�µ�������ָ�������ӿ�
	//ע�������ǸĵĶ������ݶ��Ƕ��ļĴ����ţ����AT��������ﲻӰ��
	
	///////////////////// lui Shifter ////////////////////////
	wire [31:0] luiRes_wire;
	assign luiRes_wire = {Instr[15:0], 16'd0};
	
	///////////////////// Branch ////////////////////////////
	
	assign branch = (`beq && RsData_wire == RtData_wire) ? 1 : 0;
	assign branch_addr32 = PC_4 + {imm32_wire[29:0], 2'b00};
	
	///////////////////// Jump /////////////////////////
	assign jump = (`j || `jal || `jr) ? 1 : 0;
	assign jump_addr32 = `j || `jal ? {PC[31:28], imm26_wire, 2'b00}:
	                     `jr ? RsData_wire : 32'h0000_3000;
	
	//////////////////// ��֧����ûд��/////////////////////
	assign RsData_wire = RData0_wire;
	assign RtData_wire = RData1_wire;
	////////////////// ID/EX��ˮ�߼Ĵ��� ////////////////////
	
	always@(posedge clk)
	begin
		if(reset)
		begin
			Rs_ID_to_EX <= 5'd0;
			Rt_ID_to_EX <= 5'd0;
			RegWriteAddr_ID_to_EX <= 5'd0;
			Shamt_ID_to_EX <= 5'd0;
			imm32_ID_to_EX <= 32'd0;
			InstrType_ID_to_EX <= `inst_sll; // Type of nop(sll)
			RsData_ID_to_EX <= 32'd0;
			RtData_ID_to_EX <= 32'd0;
			luiRes_ID_to_EX <= 32'd0;
			PC_ID_to_EX <= 32'h0000_3000;
		end
		else
		begin
			Rs_ID_to_EX <= Rs_wire;
			Rt_ID_to_EX <= Rt_wire;
			RegWriteAddr_ID_to_EX <= WAddr_wire; //��ǰָ����ʵ��д���ַ
			Shamt_ID_to_EX <= Shamt_wire;
			imm32_ID_to_EX <= imm32_wire;
			InstrType_ID_to_EX <= InstrType;
			RsData_ID_to_EX <= RsData_wire;
			RtData_ID_to_EX <= RtData_wire;
			luiRes_ID_to_EX <= luiRes_wire;
			PC_ID_to_EX <= PC;
		end
	end
	
endmodule
